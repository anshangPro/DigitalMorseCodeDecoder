`timescale 1ns / 1ps

module keyBoard(
input clk,
input rst,
input [3:0] row,
output reg [3:0] col,
output reg [3:0] key
    );

endmodule
