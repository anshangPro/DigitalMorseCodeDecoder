`timescale 1ns / 1ps

module encoder(
input en,
input clk,
input rst,
input [3:0] key,
input encode_button,
output [7:0] seg_en,
output [7:0] seg_out
    );

endmodule
