`timescale 1ns / 1ps

module mode_switch(
    input sw,
    output reg decoder_en,
    output reg encoder_en
);
   

decoder();
encoder();
endmodule
